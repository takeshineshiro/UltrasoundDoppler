`timescale 1ns/10ps

module tbslave;
    reg rstb = 1'b0;
    reg ten = 1'b0;
    reg [15:0] tdata = 16'h0000;
    reg mlb = 1'b0;
    reg ss = 1'b0;
    reg sck = 1'b0;
    reg sdin = 1'b0;
    wire sdout;
    wire done;
    wire [15:0] rdata;


    SPI_slave UUT (
        .rstb(rstb),
        .ten(ten),
        .tdata(tdata),
        .sck(sck),
        .mosi(sdin),
        .miso(sdout),
        .done(done),
        .rdata(rdata));

    initial begin
        // -------------  Current Time:  100ns
        #100;
        ss = 1'b1;
        sck = 1'b1;
        sdin = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  120ns
        #20;
        rstb = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  140ns
        #20;
        ten = 1'b1;
        mlb = 1'b1;
        tdata = 16'hAAAA;
        // -------------------------------------
        // -------------  Current Time:  160ns
        #20;
        ss = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  180ns
        #20;
        sck = 1'b0;
        sdin = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  200ns
        #20;
        sck = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  220ns
        #20;
        sck = 1'b0;
        sdin = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  240ns
        #20;
        sck = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  260ns
        #20;
        sck = 1'b0;
        sdin = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  280ns
        #20;
        sck = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  300ns
        #20;
        sck = 1'b0;
        sdin = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  320ns
        #20;
        sck = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  340ns
        #20;
        sck = 1'b0;
        sdin = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  360ns
        #20;
        sck = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  380ns
        #20;
        sck = 1'b0;
        sdin = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  400ns
        #20;
        sck = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  420ns
        #20;
        sck = 1'b0;
        sdin = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  440ns
        #20;
        sck = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  460ns
        #20;
        sck = 1'b0;
        sdin = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  480ns
        #20;
        sck = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  500ns
        #20;
        ss = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  520ns
        #20;
        ten = 1'b0;

		
		#200  ten = 1'b1;        mlb = 1'b0;         tdata = 16'hAFAF;
        #20        ss = 1'b0;
        #20       sck = 1'b0;
        sdin = 1'b0;
        #20        sck = 1'b1;
        #20        sck = 1'b0;
        sdin = 1'b1;
        #20        sck = 1'b1;

        #20        sck = 1'b0;
        sdin = 1'b0;
        #20        sck = 1'b1;
        #20        sck = 1'b0;
        sdin = 1'b1;
        #20        sck = 1'b1;
        #20        sck = 1'b0;
        sdin = 1'b0;
        #20        sck = 1'b1;
        #20        sck = 1'b0;
        sdin = 1'b1;
        #20        sck = 1'b1;
        #20        sck = 1'b0;
        sdin = 1'b0;
        #20        sck = 1'b1;
        #20        sck = 1'b0;
        sdin = 1'b1;
        #20        sck = 1'b1;
        #20         ss = 1'b1;
        #20         ten = 1'b0;
		#100;

	end

endmodule

